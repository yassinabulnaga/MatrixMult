// Simple DMA Controller for Matrix Transfer
// Supports: DDR -> BRAM (load) and BRAM -> DDR (store)

module dma_controller #(
    parameter int N = 16
)(
    input  logic        clk,
    input  logic        rst,
    
    // Control interface
    input  logic        start_load_a,      // Load matrix A from DDR
    input  logic        start_load_b,      // Load matrix B from DDR
    input  logic        start_store_c,     // Store matrix C to DDR
    input  logic [31:0] addr_a,            // DDR address for matrix A
    input  logic [31:0] addr_b,            // DDR address for matrix B
    input  logic [31:0] addr_c,            // DDR address for matrix C
    output logic        done,
    output logic        busy,
    
    // Avalon-MM Master to DDR (simplified)
    output logic [31:0] avm_address,
    output logic        avm_read,
    output logic        avm_write,
    output logic [31:0] avm_writedata,
    input  logic [31:0] avm_readdata,
    input  logic        avm_readdatavalid,
    input  logic        avm_waitrequest,
    output logic [3:0]  avm_byteenable,
    
    // BRAM A interface (16 banks, 8-bit each)
    output logic [15:0][7:0] bram_a_addr,
    output logic [15:0][7:0] bram_a_wdata,
    output logic [15:0]      bram_a_wren,
    
    // BRAM B interface (16 banks, 8-bit each)
    output logic [15:0][7:0] bram_b_addr,
    output logic [15:0][7:0] bram_b_wdata,
    output logic [15:0]      bram_b_wren,
    
    // BRAM C interface (16 banks, 32-bit each)
    output logic [15:0][7:0]  bram_c_addr,
    input  logic [15:0][31:0] bram_c_rdata
);

    typedef enum logic [2:0] {
        IDLE,
        LOAD_A,
        LOAD_B,
        STORE_C,
        DONE
    } state_t;
    
    state_t state_d, state_q;
    
    logic [31:0] base_addr_d, base_addr_q;
    logic [7:0]  row_cnt_d, row_cnt_q;
    logic [3:0]  col_cnt_d, col_cnt_q;
    logic        read_issued_d, read_issued_q;
    
    always_ff @(posedge clk or negedge rst) begin
        if (!rst) begin
            state_q <= IDLE;
            base_addr_q <= '0;
            row_cnt_q <= '0;
            col_cnt_q <= '0;
            read_issued_q <= 1'b0;
        end else begin
            state_q <= state_d;
            base_addr_q <= base_addr_d;
            row_cnt_q <= row_cnt_d;
            col_cnt_q <= col_cnt_d;
            read_issued_q <= read_issued_d;
        end
    end
    
    always_comb begin
        // Defaults
        state_d = state_q;
        base_addr_d = base_addr_q;
        row_cnt_d = row_cnt_q;
        col_cnt_d = col_cnt_q;
        read_issued_d = read_issued_q;
        
        avm_address = '0;
        avm_read = 1'b0;
        avm_write = 1'b0;
        avm_writedata = '0;
        avm_byteenable = 4'hF;
        
        bram_a_addr = '0;
        bram_a_wdata = '0;
        bram_a_wren = '0;
        bram_b_addr = '0;
        bram_b_wdata = '0;
        bram_b_wren = '0;
        bram_c_addr = '0;
        
        done = 1'b0;
        busy = (state_q != IDLE);
        
        case (state_q)
            IDLE: begin
                if (start_load_a) begin
                    state_d = LOAD_A;
                    base_addr_d = addr_a;
                    row_cnt_d = '0;
                    col_cnt_d = '0;
                    read_issued_d = 1'b0;
                end else if (start_load_b) begin
                    state_d = LOAD_B;
                    base_addr_d = addr_b;
                    row_cnt_d = '0;
                    col_cnt_d = '0;
                    read_issued_d = 1'b0;
                end else if (start_store_c) begin
                    state_d = STORE_C;
                    base_addr_d = addr_c;
                    row_cnt_d = '0;
                    col_cnt_d = '0;
                end
            end
            
            LOAD_A: begin
                // Issue read only if we haven't issued one yet
                if (!read_issued_q) begin
                    avm_address = base_addr_q + (row_cnt_q * N + col_cnt_q * 4);
                    avm_read = 1'b1;
                    if (!avm_waitrequest) begin
                        read_issued_d = 1'b1;
                    end
                end
                
                // When data is valid, write to BRAM
                if (avm_readdatavalid) begin
                    // Write 4 consecutive bytes to 4 consecutive banks
                    for (int i = 0; i < 4; i++) begin
                        bram_a_addr[col_cnt_q*4 + i] = row_cnt_q;
                        bram_a_wdata[col_cnt_q*4 + i] = avm_readdata[i*8 +: 8];
                        bram_a_wren[col_cnt_q*4 + i] = 1'b1;
                    end
                    
                    read_issued_d = 1'b0;  // Ready for next read
                    col_cnt_d = col_cnt_q + 1;
                    
                    if (col_cnt_q == 3) begin  // 4 reads (0,1,2,3) * 4 bytes = 16 bytes per row
                        col_cnt_d = '0;
                        if (row_cnt_q == N-1) begin
                            state_d = DONE;
                        end else begin
                            row_cnt_d = row_cnt_q + 1;
                        end
                    end
                end
            end
            
            LOAD_B: begin
                // Issue read only if we haven't issued one yet
                if (!read_issued_q) begin
                    avm_address = base_addr_q + (row_cnt_q * N + col_cnt_q * 4);
                    avm_read = 1'b1;
                    if (!avm_waitrequest) begin
                        read_issued_d = 1'b1;
                    end
                end
                
                if (avm_readdatavalid) begin
                    for (int i = 0; i < 4; i++) begin
                        bram_b_addr[col_cnt_q*4 + i] = row_cnt_q;
                        bram_b_wdata[col_cnt_q*4 + i] = avm_readdata[i*8 +: 8];
                        bram_b_wren[col_cnt_q*4 + i] = 1'b1;
                    end
                    
                    read_issued_d = 1'b0;
                    col_cnt_d = col_cnt_q + 1;
                    
                    if (col_cnt_q == 3) begin
                        col_cnt_d = '0;
                        if (row_cnt_q == N-1) begin
                            state_d = DONE;
                        end else begin
                            row_cnt_d = row_cnt_q + 1;
                        end
                    end
                end
            end
            
            STORE_C: begin
                // Read from BRAM C and write to DDR
                // Read 1 element (32-bit) at a time
                for (int i = 0; i < 16; i++) begin
                    bram_c_addr[i] = row_cnt_q;
                end
                
                // Write current column's data to DDR
                avm_address = base_addr_q + (row_cnt_q * N + col_cnt_q) * 4;  // 4 bytes per int32
                avm_write = 1'b1;
                avm_writedata = bram_c_rdata[col_cnt_q];
                
                if (!avm_waitrequest) begin
                    col_cnt_d = col_cnt_q + 1;
                    if (col_cnt_q == N-1) begin
                        col_cnt_d = '0;
                        if (row_cnt_q == N-1) begin
                            state_d = DONE;
                        end else begin
                            row_cnt_d = row_cnt_q + 1;
                        end
                    end
                end
            end
            
            DONE: begin
                done = 1'b1;
                state_d = IDLE;
            end
        endcase
    end

endmodule