// Main State Machine - Orchestrates DMA and Matrix Multiplication
// Flow: Load A -> Load B -> Compute -> Store C

module matmul_fsm #(
    parameter int N = 16
)(
    input  logic        clk,
    input  logic        rst,
    
    // Control from CPU
    input  logic        start,             // Start complete operation
    input  logic [31:0] ddr_addr_a,        // DDR address for matrix A
    input  logic [31:0] ddr_addr_b,        // DDR address for matrix B  
    input  logic [31:0] ddr_addr_c,        // DDR address for matrix C
    output logic        complete,          // Operation complete
    output logic        busy,
    
    // DMA control
    output logic        dma_start_load_a,
    output logic        dma_start_load_b,
    output logic        dma_start_store_c,
    output logic [31:0] dma_addr_a,
    output logic [31:0] dma_addr_b,
    output logic [31:0] dma_addr_c,
    input  logic        dma_done,
    input  logic        dma_busy,
    
    // Compute control
    output logic        compute_start,
    input  logic        compute_done
);

    typedef enum logic [3:0] {
        IDLE,
        LOAD_A,
        WAIT_A,
        LOAD_B,
        WAIT_B,
        COMPUTE,
        WAIT_COMPUTE,
        STORE_C,
        WAIT_STORE,
        COMPLETE
    } state_t;
    
    state_t state_d, state_q;
    
    always_ff @(posedge clk or negedge rst) begin
        if (!rst) begin
            state_q <= IDLE;
        end else begin
            state_q <= state_d;
        end
    end
    
    always_comb begin
        // Defaults
        state_d = state_q;
        
        dma_start_load_a = 1'b0;
        dma_start_load_b = 1'b0;
        dma_start_store_c = 1'b0;
        dma_addr_a = ddr_addr_a;
        dma_addr_b = ddr_addr_b;
        dma_addr_c = ddr_addr_c;
        
        compute_start = 1'b0;
        
        complete = 1'b0;
        busy = (state_q != IDLE);
        
        case (state_q)
            IDLE: begin
                if (start) begin
                    state_d = LOAD_A;
                end
            end
            
            LOAD_A: begin
                dma_start_load_a = 1'b1;
                state_d = WAIT_A;
            end
            
            WAIT_A: begin
                if (dma_done) begin
                    state_d = LOAD_B;
                end
            end
            
            LOAD_B: begin
                dma_start_load_b = 1'b1;
                state_d = WAIT_B;
            end
            
            WAIT_B: begin
                if (dma_done) begin
                    state_d = COMPUTE;
                end
            end
            
            COMPUTE: begin
                compute_start = 1'b1;
                state_d = WAIT_COMPUTE;
            end
            
            WAIT_COMPUTE: begin
                if (compute_done) begin
                    state_d = STORE_C;
                end
            end
            
            STORE_C: begin
                dma_start_store_c = 1'b1;
                state_d = WAIT_STORE;
            end
            
            WAIT_STORE: begin
                if (dma_done) begin
                    state_d = COMPLETE;
                end
            end
            
            COMPLETE: begin
                complete = 1'b1;
                state_d = IDLE;
            end
        endcase
    end

endmodule