`timescale 1ns/1ps

module tb_fifo_wrapper;

  // Parameters
  localparam int W = 16;        // Data width for matrix elements
  localparam int LGFLEN = 7;    // 2^7 = 128 depth FIFO
  localparam int DEPTH = 1 << LGFLEN;
  
  // DUT signals
  logic clk, rst_n;
  logic [W-1:0] s_data;         // Slave (input) interface
  logic         s_valid;
  logic         s_ready;
  logic [W-1:0] m_data;         // Master (output) interface  
  logic         m_valid;
  logic         m_ready;
  
  // Test variables
  int i, j;
  int errors = 0;
  logic [W-1:0] test_data[$];   // Queue for checking
  logic [W-1:0] received_data;
  int write_count, read_count;
int total_elems;

  
  // Clock generation - 100MHz
  initial clk = 0;
  always #5 clk = ~clk;
  
  // DUT instantiation
  fifo_wrapper #(
    .W(W),
    .LGFLEN(LGFLEN)
  ) DUT (
    .clk(clk),
    .rst_n(rst_n),
    .s_data(s_data),
    .s_valid(s_valid),
    .s_ready(s_ready),
    .m_data(m_data),
    .m_valid(m_valid),
    .m_ready(m_ready)
  );
  
  // Reset task
  task reset_dut();
    rst_n = 0;
    s_valid = 0;
    m_ready = 0;
    s_data = '0;
    @(posedge clk);
    @(posedge clk);
    rst_n = 1;
    @(posedge clk);
  endtask
  
  // Write task - simulates drainer pushing data
  task write_data(input logic [W-1:0] data);
    s_data = data;
    s_valid = 1;
    @(posedge clk);
    while (!s_ready) @(posedge clk);  // Wait if FIFO full
    s_valid = 0;
  endtask
  
task read_data(output logic [W-1:0] data);
  m_ready = 1;

  // Wait until data is valid (with ready already high),
  // so handshake (m_valid && m_ready) happens on this cycle.
  @(posedge clk);
  while (!m_valid) @(posedge clk);

  data    = m_data;  // capture the word from the handshake cycle
  m_ready = 0;
endtask

  
  // Continuous write task (with backpressure handling)
  task automatic continuous_write(input int count, input int start_val);
    automatic int k;
    for (k = 0; k < count; k++) begin
      s_data = start_val + k;
      s_valid = 1;
      @(posedge clk);
      if (s_ready) begin
        test_data.push_back(start_val + k);
        write_count++;
      end else begin
        k--;  // Retry if not ready
      end
    end
    s_valid = 0;
  endtask
  
  // Continuous read task (with flow control)
  task automatic continuous_read(input int count);
    automatic int k;
    for (k = 0; k < count; k++) begin
      m_ready = 1;
      @(posedge clk);
      if (m_valid) begin
        received_data = m_data;
        if (test_data.size() > 0) begin
          automatic logic [W-1:0] expected_val = test_data.pop_front();
          if (received_data !== expected_val) begin
            $error("[FAIL] Data mismatch at read %0d: got %h, expected %h",
                   k, received_data, expected_val);
            errors++;
          end
        end
        read_count++;
      end else begin
        k--;  // Retry if no valid data
      end
    end
    m_ready = 0;
  endtask
  
  // Main test
  initial begin
    $display("=== FIFO Wrapper Testbench for Matrix Multiplier ===");
    $display("FIFO Depth: %0d, Data Width: %0d bits", DEPTH, W);
    
    // Initialize
    reset_dut();
    test_data.delete();
    write_count = 0;
    read_count = 0;
    
    //==================================================================
    // Test 1: Basic write and read
    //==================================================================
    $display("\n[Test 1] Basic write and read");
    
    // Write 10 values
    for (i = 0; i < 10; i++) begin
      write_data(16'h1000 + i);
      test_data.push_back(16'h1000 + i);
    end
    
    // Read 10 values
    for (i = 0; i < 10; i++) begin
      automatic logic [W-1:0] expected_val = test_data.pop_front();
      read_data(received_data);
      if (received_data !== expected_val) begin
        $error("[FAIL] Test 1: Data mismatch at %0d", i);
        errors++;
      end
    end
    
    $display("[PASS] Test 1: Basic write/read OK");
$display("Time = %0t ns", $time);

    
    //==================================================================
// Test 2: Fill FIFO completely (test full condition)
//==================================================================
$display("\n[Test 2] Fill FIFO to full");
reset_dut();
test_data.delete();

i = 0;

// Drive until we get DEPTH *accepted* writes
while (i < DEPTH) begin
  s_valid = 1;
  s_data  = i[W-1:0];

  @(posedge clk);

  if (s_ready) begin
    // Handshake happened this cycle: s_valid && s_ready
    test_data.push_back(i[W-1:0]);
    i++;
  end
  // else: FIFO is full this cycle; keep s_valid high and retry
end

// Stop driving valid
s_valid = 0;

// Give FIFO one clock to update full flag
@(posedge clk);

// Now s_ready must be low if FIFO is full
if (s_ready) begin
  $error("[FAIL] Test 2: s_ready should be 0 when FIFO is full (accepted %0d)", test_data.size());
  errors++;
end else begin
  $display("[PASS] Test 2: FIFO full detection works (accepted %0d entries)", test_data.size());
$display("Time = %0t ns", $time);

end

    
    //==================================================================
    // Test 3: Empty FIFO completely (test empty condition)  
    //==================================================================
    $display("\n[Test 3] Empty FIFO completely");
    
    // Read all data
    while (test_data.size() > 0) begin
      automatic logic [W-1:0] expected_val = test_data.pop_front();
      read_data(received_data);
      if (received_data !== expected_val) begin
        $error("[FAIL] Test 3: Data mismatch");
        errors++;
      end
    end
@(posedge clk);  // allow empty/m_valid to update

    
    // Verify m_valid deasserted when empty
    if (m_valid) begin
      $error("[FAIL] Test 3: m_valid should be 0 when FIFO is empty");
$display("Time = %0t ns", $time);

      errors++;
    end else begin
      $display("[PASS] Test 3: FIFO empty detection works");
    end
    
    //==================================================================
    // Test 4: Simultaneous read/write (streaming)
    //==================================================================
    $display("\n[Test 4] Simultaneous read/write (matrix data streaming)");
    reset_dut();
    test_data.delete();
    write_count = 0;
    read_count = 0;
    
    // Simulate continuous data flow from drainer to packer
    fork
      // Writer thread (simulates drainer)
      begin
        continuous_write(256, 16'hA000);
      end
      
      // Reader thread (simulates packer)
      begin
        #50;  // Small delay to let some data accumulate
        continuous_read(256);
      end
    join
    
    $display("[INFO] Test 4: Wrote %0d, Read %0d", write_count, read_count);
    if (write_count == 256 && read_count == 256 && errors == 0) begin
      $display("[PASS] Test 4: Streaming operation successful");
    end else begin
      $error("[FAIL] Test 4: Streaming mismatch");
      errors++;
    end
    
    //==================================================================
    // Test 5: Burst write with slow read (backpressure test)
    //==================================================================
    $display("\n[Test 5] Burst write with slow read (backpressure)");
    reset_dut();
    test_data.delete();
    
    // Write burst of data
    fork
      begin
        for (i = 0; i < 200; i++) begin
          s_data = 16'hB000 | i[W-1:0];
          s_valid = 1;
          @(posedge clk);
          if (s_ready) test_data.push_back(16'hB000 | i[W-1:0]);
          else i--;  // Retry
        end
        s_valid = 0;
      end
      
      // Slow reader
      begin
        automatic int k;
        repeat(10) @(posedge clk);
        for (k = 0; k < 200; k++) begin
          m_ready = 1;
          @(posedge clk);
          if (m_valid) begin
            automatic logic [W-1:0] expected_val;
            received_data = m_data;
            expected_val = test_data.pop_front();
            if (received_data !== expected_val) begin
              $error("[FAIL] Test 5: Data mismatch at %0d", k);
              errors++;
            end
          end else begin
            k--;
          end
          m_ready = 0;
          repeat(2) @(posedge clk);  // Slow read rate
        end
      end
    join
    
    $display("[PASS] Test 5: Backpressure handling OK");
    
//==================================================================
// Test 6: Matrix data pattern (16x16 matrix)
//==================================================================
$display("\n[Test 6] Matrix data pattern (16x16 matrix)");
reset_dut();
test_data.delete();      // not used here, but okay to clear
write_count  = 0;
read_count   = 0;
total_elems  = 16*16;

// We stream 256 elements through the 128-deep FIFO using
// concurrent writer and reader. At no point do we require
// more than DEPTH entries in-flight.
fork
  // ---------------- Writer thread ----------------
  begin
    int r, c;
    logic [W-1:0] val;

    for (r = 0; r < 16; r = r + 1) begin
      for (c = 0; c < 16; c = c + 1) begin
        val     = (r << 8) | c;
        s_data  = val;
        s_valid = 1;

        // Wait for handshake s_valid && s_ready
        @(posedge clk);
        while (!s_ready) @(posedge clk);

        write_count++;

        s_valid = 0;
        // optional small gap; can be removed if you want max throughput
        // @(posedge clk);
      end
    end

    s_valid = 0;
  end

  // ---------------- Reader thread ----------------
  begin
    int k;
    logic [W-1:0] got, exp;

    // Let writer start
    @(posedge clk);

    for (k = 0; k < total_elems; k = k + 1) begin
      m_ready = 1;

      // Wait for handshake m_valid && m_ready
      @(posedge clk);
      while (!m_valid) @(posedge clk);

      got = m_data;

      // Reconstruct expected [row][col] for index k
      exp = ((k / 16) << 8) | (k % 16);

      if (got !== exp) begin
        $error("[FAIL] Test 6: mismatch at index %0d: got %h, expected %h",
               k, got, exp);
        errors++;
      end

      read_count++;
    end

    m_ready = 0;
  end
join

// Let empty/m_valid settle
@(posedge clk);

$display("[INFO] Test 6: Wrote %0d, Read %0d", write_count, read_count);
if (write_count == total_elems && read_count == total_elems && errors == 0 && !m_valid) begin
  $display("[PASS] Test 6: Matrix streaming pattern OK");
end else begin
  $error("[FAIL] Test 6: Matrix streaming / count mismatch");
end


    
    //==================================================================
    // Test 7: Reset during operation
    //==================================================================
    $display("\n[Test 7] Reset during operation");
    
    // Fill partially
    for (i = 0; i < 50; i++) begin
      write_data(16'hCC00 + i);
    end
    
    // Reset while data is in FIFO
    reset_dut();
    
    // Check that FIFO is empty after reset
    if (m_valid) begin
      $error("[FAIL] Test 7: FIFO should be empty after reset");
      errors++;
    end else begin
      $display("[PASS] Test 7: Reset clears FIFO properly");
    end
    
    //==================================================================
    // Test 8: Single-cycle write/read transitions
    //==================================================================
    $display("\n[Test 8] Single-cycle transitions");
    reset_dut();
    
    // Rapid write-read-write-read pattern
    for (i = 0; i < 20; i++) begin
      // Write
      s_data = 16'hDD00 + i;
      s_valid = 1;
      m_ready = 0;
      @(posedge clk);
      s_valid = 0;
      
      // Read
      m_ready = 1;
      @(posedge clk);
      if (m_valid && m_data !== (16'hDD00 + i)) begin
        $error("[FAIL] Test 8: Fast transition mismatch at %0d", i);
        errors++;
      end
      m_ready = 0;
      @(posedge clk);
    end
    
    $display("[PASS] Test 8: Single-cycle transitions OK");
    
    //==================================================================
    // Final Report
    //==================================================================
    $display("\n============================================================");
    if (errors == 0) begin
      $display("ALL TESTS PASSED!");
    end else begin
      $display("TESTS FAILED with %0d errors", errors);
    end
    $display("============================================================");
    
    $finish;
  end
  
  // Timeout watchdog
  initial begin
    #100000;  // 100us timeout
    $error("Test timeout!");
`    $finish;
  end
  
  // Optional: Monitor FIFO fill level (commented out to reduce verbosity)
  /*
  always @(posedge clk) begin
    if (rst_n && (s_valid || m_ready)) begin
      $display("[%0t] s_valid=%b s_ready=%b | m_valid=%b m_ready=%b | data=%h", 
               $time, s_valid, s_ready, m_valid, m_ready, 
               s_valid ? s_data : m_data);
    end
  end
  */

endmodule