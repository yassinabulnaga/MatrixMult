module dp_bram #(
    parameter int W           = 128,
    parameter int DEPTH       = 1024,
    parameter bit USE_BYTE_EN = 1,
    parameter int AW          = (DEPTH <= 1) ? 1 : $clog2(DEPTH),
    // 0 = WRITE_FIRST, 1 = READ_FIRST, 2 = NO_CHANGE
    parameter int RDW_MODE    = 2
)(
    input  logic              clk,
    input  logic              rst_n,

    // Port A
    input  logic              a_en,
    input  logic [AW-1:0]     a_addr,
    input  logic [W-1:0]      a_din,
    input  logic              a_we,
    input  logic [W/8-1:0]    a_be,
    output logic [W-1:0]      a_dout,

    // Port B
    input  logic              b_en,
    input  logic [AW-1:0]     b_addr,
    input  logic [W-1:0]      b_din,
    input  logic              b_we,
    input  logic [W/8-1:0]    b_be,
    output logic [W-1:0]      b_dout
);

  (* ramstyle = "M10K, no_rw_check" *)
  logic [W-1:0] mem [0:DEPTH-1];

  logic [W-1:0] a_q, b_q;

  // Sanity checks
  initial begin
    if (USE_BYTE_EN && (W % 8) != 0)
      $fatal(1, "dp_bram: W must be multiple of 8 when USE_BYTE_EN=1");
    if (RDW_MODE < 0 || RDW_MODE > 2)
      $fatal(1, "dp_bram: RDW_MODE must be 0/1/2");
  end

  // Byte-enable helper
  function automatic [W-1:0] mask_write(
      input [W-1:0]    din,
      input [W-1:0]    prev,
      input [W/8-1:0]  be
  );
    if (!USE_BYTE_EN) begin
      return din;
    end else begin
      automatic logic [W-1:0] res;
      int i;
      for (i = 0; i < W/8; i++) begin
        res[i*8 +: 8] = be[i] ? din[i*8 +: 8] : prev[i*8 +: 8];
      end
      return res;
    end
  endfunction

  // Port A
  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      a_q <= '0;
    end else if (a_en) begin
      automatic logic [W-1:0] prev;
      automatic logic [W-1:0] wdata;

      prev  = mem[a_addr];
      wdata = mask_write(a_din, prev, a_be);

      if (a_we)
        mem[a_addr] <= wdata;

      unique case (RDW_MODE)
        0: a_q <= a_we ? wdata : prev;     // WRITE_FIRST
        1: a_q <= prev;                    // READ_FIRST (old data)
        2: a_q <= a_we ? a_q : prev;       // NO_CHANGE on write
        default: a_q <= prev;
      endcase
    end
  end

  // Port B
  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      b_q <= '0;
    end else if (b_en) begin
      automatic logic [W-1:0] prev;
      automatic logic [W-1:0] wdata;

      prev  = mem[b_addr];
      wdata = mask_write(b_din, prev, b_be);

      if (b_we)
        mem[b_addr] <= wdata;

      unique case (RDW_MODE)
        0: b_q <= b_we ? wdata : prev;     // WRITE_FIRST
        1: b_q <= prev;                    // READ_FIRST
        2: b_q <= b_we ? b_q : prev;       // NO_CHANGE
        default: b_q <= prev;
      endcase
    end
  end

  // Output pipeline stage (kept for timing / M10K style)
  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      a_dout <= '0;
      b_dout <= '0;
    end else begin
      a_dout <= a_q;
      b_dout <= b_q;
    end
  end

endmodule

